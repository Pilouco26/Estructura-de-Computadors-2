//: version "1.8.7"

module UC(MemToReg, MemWrite, MemRead, Branch, RegDst, RegWrite, Jump, AluSrc, AluOp, op);
//: interface  /sz:(238, 91) /bd:[ Li0>op[5:0](36/91) To0<Jump(223/238) Lo0<RegDst(22/91) Bo0<RegWrite(176/238) Ro0<Branch(14/91) Ro1<MemRead(29/91) Ro2<MemToReg(39/91) Ro3<AluOp[1:0](53/91) Ro4<MemWrite(65/91) Ro5<AluSrc(77/91) ]
output Branch;    //: /sn:0 {0}(709,326)(709,303)(621,303){1}
//: {2}(619,301)(619,274){3}
//: {4}(621,272)(671,272)(671,335){5}
//: {6}(669,337)(648,337)(648,361){7}
//: {8}(671,339)(671,393){9}
//: {10}(619,270)(619,204){11}
//: {12}(619,305)(619,314){13}
output MemWrite;    //: /sn:0 {0}(937,301)(937,244){1}
output AluSrc;    //: /sn:0 /dp:1 {0}(692,274)(692,254)(699,254){1}
//: {2}(703,254)(714,254)(714,268){3}
//: {4}(716,270)(777,270)(777,331){5}
//: {6}(714,272)(714,326){7}
//: {8}(701,252)(701,204){9}
//: {10}(701,256)(701,281)(733,281)(733,362){11}
output RegDst;    //: /sn:0 {0}(661,393)(661,369)(707,369){1}
//: {2}(709,367)(709,347){3}
//: {4}(709,371)(709,387){5}
output RegWrite;    //: /sn:0 {0}(619,405)(619,370){1}
output MemRead;    //: /sn:0 /dp:1 {0}(780,388)(780,352){1}
output [1:0] AluOp;    //: /sn:0 /dp:1 {0}(666,399)(666,432){1}
output MemToReg;    //: /sn:0 {0}(888,303)(888,265){1}
//: {2}(888,261)(888,204){3}
//: {4}(886,263)(820,263)(820,280){5}
input [5:0] op;    //: /sn:0 /dp:1 {0}(557,200)(601,200){1}
//: {2}(602,200)(618,200){3}
//: {4}(619,200)(638,200){5}
//: {6}(639,200)(655,200){7}
//: {8}(656,200)(680,200)(680,200)(700,200){9}
//: {10}(701,200)(830,200){11}
//: {12}(831,200)(887,200){13}
//: {14}(888,200)(912,200)(912,240)(936,240){15}
//: {16}(937,240)(1104,240){17}
output Jump;    //: /sn:0 {0}(829,377)(829,331){1}
wire w6;    //: /sn:0 /dp:1 {0}(619,354)(619,335){1}
wire w7;    //: /sn:0 /dp:1 {0}(614,314)(614,275)(642,275)(642,265){1}
wire w4;    //: /sn:0 {0}(820,296)(820,308)(826,308)(826,310){1}
wire w3;    //: /sn:0 /dp:1 {0}(656,215)(656,195){1}
wire w0;    //: /sn:0 /dp:1 {0}(624,314)(624,313)(689,313)(689,295){1}
wire w1;    //: /sn:0 /dp:1 {0}(639,244)(639,204){1}
wire w11;    //: /sn:0 {0}(656,231)(656,241)(644,241)(644,244){1}
wire w2;    //: /sn:0 /dp:1 {0}(831,310)(831,204){1}
wire Jump1;    //: /sn:0 {0}(687,274)(687,263){1}
//: {2}(689,261)(782,261)(782,269){3}
//: {4}(685,261)(604,261){5}
//: {6}(602,259)(602,204){7}
//: {8}(602,263)(602,279)(704,279)(704,326){9}
wire w5;    //: /sn:0 /dp:1 {0}(782,331)(782,285){1}
//: enddecls

  //: output g4 (MemToReg) @(888,300) /sn:0 /R:3 /w:[ 0 ]
  //: output g8 (MemWrite) @(937,298) /sn:0 /R:3 /w:[ 0 ]
  //: output g3 (MemRead) @(780,385) /sn:0 /R:3 /w:[ 0 ]
  tran g16(.Z(AluSrc), .I(op[5]));   //: @(701,198) /sn:0 /R:1 /w:[ 9 9 10 ] /ss:1
  tran g26(.Z(w2), .I(op[1]));   //: @(831,198) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  not g17 (.I(w6), .Z(RegWrite));   //: @(619,360) /sn:0 /R:3 /w:[ 0 1 ]
  //: output g2 (Branch) @(648,358) /sn:0 /R:3 /w:[ 7 ]
  concat g23 (.I0(Branch), .I1(RegDst), .Z(AluOp));   //: @(666,398) /sn:0 /R:3 /w:[ 9 0 0 ] /dr:1
  //: joint g30 (Jump1) @(602, 261) /w:[ 5 6 -1 8 ]
  //: output g1 (RegDst) @(709,384) /sn:0 /R:3 /w:[ 5 ]
  //: joint g24 (Branch) @(619, 272) /w:[ 4 10 -1 3 ]
  not g29 (.I(Jump1), .Z(w5));   //: @(782,275) /sn:0 /R:3 /w:[ 3 1 ]
  nor g18 (.I0(AluSrc), .I1(Branch), .I2(Jump1), .Z(RegDst));   //: @(709,337) /sn:0 /R:3 /w:[ 7 0 9 3 ]
  //: output g10 (RegWrite) @(619,402) /sn:0 /R:3 /w:[ 0 ]
  //: joint g25 (Branch) @(671, 337) /w:[ -1 5 6 8 ]
  //: output g6 (Jump) @(829,374) /sn:0 /R:3 /w:[ 0 ]
  //: joint g35 (Jump1) @(687, 261) /w:[ 2 -1 4 1 ]
  and g7 (.I0(w4), .I1(w2), .Z(Jump));   //: @(829,321) /sn:0 /R:3 /w:[ 1 0 1 ]
  //: output g9 (AluSrc) @(733,359) /sn:0 /R:3 /w:[ 11 ]
  not g31 (.I(MemToReg), .Z(w4));   //: @(820,286) /sn:0 /R:3 /w:[ 5 0 ]
  //: joint g22 (RegDst) @(709, 369) /w:[ -1 2 1 4 ]
  tran g36(.Z(w3), .I(op[0]));   //: @(656,198) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:0
  tran g33(.Z(MemToReg), .I(op[5]));   //: @(888,198) /sn:0 /R:1 /w:[ 3 13 14 ] /ss:1
  tran g12(.Z(Jump1), .I(op[3]));   //: @(602,198) /sn:0 /R:1 /w:[ 7 1 2 ] /ss:1
  //: joint g34 (MemToReg) @(888, 263) /w:[ -1 2 4 1 ]
  //: joint g28 (AluSrc) @(714, 270) /w:[ 4 3 -1 6 ]
  //: output g5 (AluOp) @(666,429) /sn:0 /R:3 /w:[ 1 ]
  or g11 (.I0(w0), .I1(Branch), .I2(w7), .Z(w6));   //: @(619,325) /sn:0 /R:3 /w:[ 0 13 0 1 ]
  and g14 (.I0(AluSrc), .I1(Jump1), .Z(w0));   //: @(689,285) /sn:0 /R:3 /w:[ 0 0 1 ]
  and g21 (.I0(w1), .I1(w11), .Z(w7));   //: @(642,255) /sn:0 /R:3 /w:[ 0 1 1 ]
  //: joint g19 (AluSrc) @(701, 254) /w:[ 2 8 1 10 ]
  //: joint g20 (Branch) @(619, 303) /w:[ 1 2 -1 12 ]
  tran g32(.Z(MemWrite), .I(op[3]));   //: @(937,238) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  //: input g0 (op) @(555,200) /sn:0 /w:[ 0 ]
  tran g15(.Z(w1), .I(op[1]));   //: @(639,198) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  and g27 (.I0(AluSrc), .I1(w5), .Z(MemRead));   //: @(780,342) /sn:0 /R:3 /w:[ 5 0 1 ]
  not g37 (.I(w3), .Z(w11));   //: @(656,221) /sn:0 /R:3 /w:[ 0 0 ]
  tran g13(.Z(Branch), .I(op[2]));   //: @(619,198) /sn:0 /R:1 /w:[ 11 3 4 ] /ss:1

endmodule

module ALU(B, A, Z, ALU_C, S);
//: interface  /sz:(72, 84) /bd:[ Li0>A[31:0](22/84) Li1>B[31:0](57/84) Bi0>ALU_C[3:0](36/72) To0<Z(48/72) Ro0<S[31:0](45/84) ]
supply0 [31:0] w7;    //: /sn:0 {0}(41,418)(41,317)(106,317){1}
input [31:0] B;    //: /sn:0 /dp:3 {0}(-358,558)(-358,464){1}
//: {2}(-356,462)(-277,462){3}
//: {4}(-358,460)(-358,349){5}
//: {6}(-356,347)(-276,347)(-276,368)(-200,368){7}
//: {8}(-358,345)(-358,289){9}
//: {10}(-356,287)(-197,287){11}
//: {12}(-358,285)(-358,273){13}
//: {14}(-356,271)(-197,271){15}
//: {16}(-358,269)(-358,245){17}
supply0 [31:0] w4;    //: /sn:0 /dp:1 {0}(106,287)(34,287)(34,289)(-37,289){1}
supply1 w0;    //: /sn:0 {0}(-202,397)(-202,422){1}
input [31:0] A;    //: /sn:0 {0}(-341,568)(-341,432){1}
//: {2}(-339,430)(-216,430){3}
//: {4}(-341,428)(-341,317){5}
//: {6}(-339,315)(-269,315)(-269,336)(-200,336){7}
//: {8}(-341,313)(-341,284){9}
//: {10}(-339,282)(-197,282){11}
//: {12}(-341,280)(-341,268){13}
//: {14}(-339,266)(-197,266){15}
//: {16}(-341,264)(-341,246){17}
output Z;    //: /sn:0 /dp:1 {0}(189,226)(189,165)(187,165)(187,160){1}
supply0 [31:0] w1;    //: /sn:0 /dp:1 {0}(106,299)(15,299)(15,304)(-54,304){1}
supply0 w8;    //: /sn:0 {0}(-186,308)(-186,328){1}
input [3:0] ALU_C;    //: /sn:0 /dp:1 {0}(122,482)(122,316){1}
supply0 [31:0] w5;    //: /sn:0 {0}(-50,296)(28,296)(28,293)(106,293){1}
output [31:0] S;    //: /sn:0 /dp:1 {0}(135,293)(187,293){1}
//: {2}(191,293)(243,293){3}
//: {4}(189,291)(189,247){5}
supply0 [30:0] w9;    //: /sn:0 {0}(-117,487)(-33,487){1}
wire w6;    //: /sn:0 {0}(-186,376)(-186,386){1}
wire [31:0] w16;    //: /sn:0 {0}(106,281)(-15,281)(-15,352)(-171,352){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(-176,285)(-36,285)(-36,275)(106,275){1}
wire [31:0] w12;    //: /sn:0 {0}(-187,446)(-97,446){1}
//: {2}(-96,446)(9,446)(9,312)(17,312)(17,305)(106,305){3}
wire [31:0] w17;    //: /sn:0 /dp:1 {0}(-27,492)(26,492)(26,311)(106,311){1}
wire w14;    //: /sn:0 {0}(-202,470)(-202,480){1}
wire w11;    //: /sn:0 {0}(-96,450)(-96,497)(-33,497){1}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(-176,269)(106,269){1}
wire [31:0] w15;    //: /sn:0 /dp:1 {0}(-261,462)(-216,462){1}
//: enddecls

  //: joint g4 (A) @(-341, 266) /w:[ 14 16 -1 13 ]
  //: joint g8 (B) @(-358, 287) /w:[ 10 12 -1 9 ]
  //: input g3 (B) @(-358,243) /sn:0 /R:3 /w:[ 17 ]
  //: supply0 g16 (w1) @(-60,304) /sn:0 /R:3 /w:[ 1 ]
  //: supply1 g26 (w0) @(-191,397) /sn:0 /w:[ 0 ]
  //: supply0 g17 (w4) @(-43,289) /sn:0 /R:3 /w:[ 1 ]
  and g2 (.I0(A), .I1(B), .Z(w2));   //: @(-186,269) /sn:0 /w:[ 15 15 0 ]
  mux g30 (.I0(w2), .I1(w3), .I2(w16), .I3(w4), .I4(w5), .I5(w1), .I6(w12), .I7(w17), .I8(w7), .S(ALU_C), .Z(S));   //: @(122,293) /sn:0 /R:1 /w:[ 1 1 0 0 1 0 3 1 1 1 0 ] /ss:0 /do:1
  //: joint g23 (S) @(189, 293) /w:[ 2 4 1 -1 ]
  //: joint g24 (B) @(-358, 462) /w:[ 2 4 -1 1 ]
  //: input g1 (A) @(-341,244) /sn:0 /R:3 /w:[ 17 ]
  //: supply0 g18 (w9) @(-123,487) /sn:0 /R:3 /w:[ 0 ]
  //: output g25 (Z) @(187,163) /sn:0 /R:1 /w:[ 1 ]
  //: joint g10 (A) @(-341, 315) /w:[ 6 8 -1 5 ]
  or g6 (.I0(A), .I1(B), .Z(w3));   //: @(-186,285) /sn:0 /w:[ 11 11 0 ]
  //: joint g7 (A) @(-341, 282) /w:[ 10 12 -1 9 ]
  add g9 (.A(B), .B(A), .S(w16), .CI(w8), .CO(w6));   //: @(-184,352) /sn:0 /R:1 /w:[ 7 7 1 1 0 ]
  nor g22 (.I0(S), .Z(Z));   //: @(189,236) /sn:0 /R:1 /w:[ 5 0 ]
  add g12 (.A(w15), .B(A), .S(w12), .CI(w0), .CO(w14));   //: @(-200,446) /sn:0 /R:1 /w:[ 1 3 0 1 0 ]
  tran g28(.Z(w11), .I(w12[31]));   //: @(-96,444) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g5 (B) @(-358, 271) /w:[ 14 16 -1 13 ]
  //: joint g11 (B) @(-358, 347) /w:[ 6 8 -1 5 ]
  //: supply0 g14 (w5) @(-56,296) /sn:0 /R:3 /w:[ 0 ]
  not g21 (.I(B), .Z(w15));   //: @(-271,462) /sn:0 /w:[ 3 0 ]
  //: supply0 g19 (w7) @(41,424) /sn:0 /w:[ 0 ]
  //: joint g20 (A) @(-341, 430) /w:[ 2 4 -1 1 ]
  //: input g0 (ALU_C) @(122,484) /sn:0 /R:1 /w:[ 0 ]
  //: output g15 (S) @(240,293) /sn:0 /w:[ 3 ]
  concat g27 (.I0(w11), .I1(w9), .Z(w17));   //: @(-28,492) /sn:0 /w:[ 1 1 0 ] /dr:0
  //: supply0 g13 (w8) @(-186,302) /sn:0 /R:2 /w:[ 0 ]

endmodule

module AC(AluCtrl, AluOp, Funct);
//: interface  /sz:(40, 40) /bd:[ ]
output [3:0] AluCtrl;    //: /sn:0 /dp:1 {0}(235,280)(235,336){1}
input [5:0] Funct;    //: /sn:0 /dp:7 {0}(389,17)(319,17){1}
//: {2}(318,17)(257,17){3}
//: {4}(256,17)(223,17){5}
//: {6}(222,17)(206,17){7}
//: {8}(205,17)(186,17){9}
//: {10}(185,17)(136,17){11}
//: {12}(135,17)(79,17){13}
supply0 w8;    //: /sn:0 {0}(250,274)(250,257){1}
input [1:0] AluOp;    //: /sn:0 {0}(80,34)(162,34){1}
//: {2}(163,34)(272,34){3}
//: {4}(273,34)(347,34){5}
//: {6}(348,34)(368,34){7}
//: {8}(369,34)(404,34){9}
wire w13;    //: /sn:0 {0}(268,112)(268,101)(257,101)(257,21){1}
wire w6;    //: /sn:0 {0}(136,21)(136,90)(108,90)(108,110){1}
wire w16;    //: /sn:0 {0}(110,131)(110,141)(145,141)(145,143){1}
wire w4;    //: /sn:0 /dp:1 {0}(230,274)(230,248)(212,248)(212,152){1}
wire w3;    //: /sn:0 {0}(273,38)(273,112){1}
wire w0;    //: /sn:0 /dp:1 {0}(298,63)(346,63){1}
//: {2}(348,61)(348,38){3}
//: {4}(348,65)(348,136)(295,136)(295,177){5}
wire w12;    //: /sn:0 /dp:1 {0}(298,58)(319,58)(319,21){1}
wire w18;    //: /sn:0 {0}(163,38)(163,113)(157,113)(157,139)(150,139)(150,143){1}
wire w10;    //: /sn:0 /dp:1 {0}(198,60)(198,42)(223,42)(223,21){1}
wire w21;    //: /sn:0 {0}(292,198)(292,217)(240,217)(240,274){1}
wire w1;    //: /sn:0 {0}(207,131)(207,115)(235,115)(235,60)(277,60){1}
wire w17;    //: /sn:0 {0}(270,133)(270,167)(290,167)(290,177){1}
wire w14;    //: /sn:0 {0}(147,164)(147,251)(220,251)(220,274){1}
wire w11;    //: /sn:0 /dp:1 {0}(196,81)(196,97)(212,97)(212,131){1}
wire w2;    //: /sn:0 /dp:1 {0}(369,69)(369,38){1}
wire w15;    //: /sn:0 {0}(193,60)(193,40)(206,40)(206,21){1}
wire w5;    //: /sn:0 {0}(186,12)(186,4)(113,4)(113,110){1}
wire w9;    //: /sn:0 {0}(369,85)(369,90)(217,90)(217,131){1}
//: enddecls

  or g8 (.I0(w9), .I1(w11), .I2(w1), .Z(w4));   //: @(212,142) /sn:0 /R:3 /w:[ 1 1 0 1 ]
  or g4 (.I0(w0), .I1(w12), .Z(w1));   //: @(287,60) /sn:0 /R:2 /w:[ 0 0 1 ]
  not g3 (.I(w2), .Z(w9));   //: @(369,75) /sn:0 /R:3 /w:[ 0 0 ]
  tran g16(.Z(w6), .I(Funct[0]));   //: @(136,15) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:1
  tran g17(.Z(w5), .I(Funct[3]));   //: @(186,15) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:0
  //: output g2 (AluCtrl) @(235,333) /sn:0 /R:3 /w:[ 1 ]
  tran g23(.Z(w18), .I(AluOp[1]));   //: @(163,32) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: input g1 (AluOp) @(78,34) /sn:0 /w:[ 0 ]
  and g18 (.I0(w18), .I1(w16), .Z(w14));   //: @(147,154) /sn:0 /R:3 /w:[ 1 1 0 ]
  tran g10(.Z(w15), .I(Funct[1]));   //: @(206,15) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  concat g6 (.I0(w14), .I1(w4), .I2(w21), .I3(w8), .Z(AluCtrl));   //: @(235,279) /sn:0 /R:3 /w:[ 1 0 1 0 0 ] /dr:0
  //: supply0 g7 (w8) @(250,251) /sn:0 /R:2 /w:[ 1 ]
  tran g9(.Z(w0), .I(AluOp[0]));   //: @(348,32) /sn:0 /R:1 /w:[ 3 5 6 ] /ss:1
  //: joint g22 (w0) @(348, 63) /w:[ -1 2 1 4 ]
  nor g12 (.I0(w10), .I1(w15), .Z(w11));   //: @(196,71) /sn:0 /R:3 /w:[ 0 0 0 ]
  tran g5(.Z(w2), .I(AluOp[1]));   //: @(369,32) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g11(.Z(w10), .I(Funct[2]));   //: @(223,15) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g14(.Z(w12), .I(Funct[1]));   //: @(319,15) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g19(.Z(w3), .I(AluOp[1]));   //: @(273,32) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g21(.Z(w13), .I(Funct[1]));   //: @(257,15) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  or g20 (.I0(w0), .I1(w17), .Z(w21));   //: @(292,188) /sn:0 /R:3 /w:[ 5 1 0 ]
  //: input g0 (Funct) @(77,17) /sn:0 /w:[ 13 ]
  or g15 (.I0(w5), .I1(w6), .Z(w16));   //: @(110,121) /sn:0 /R:3 /w:[ 1 1 0 ]
  and g13 (.I0(w3), .I1(w13), .Z(w17));   //: @(270,123) /sn:0 /R:3 /w:[ 1 0 0 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Li0>Read1[4:0](32/182) Li1>Read2[4:0](72/182) Li2>Write[4:0](108/182) Li3>WriteData[31:0](148/182) Bi0>clk(108/147) Bi1>RegWrite(40/147) Ro0<Data1[31:0](47/182) Ro1<Data2[31:0](139/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input RegWrite;    //: /sn:0 {0}(-237,263)(-172,263){1}
//: {2}(-168,263)(-71,263){3}
//: {4}(-67,263)(171,263){5}
//: {6}(175,263)(370,263){7}
//: {8}(374,263)(552,263)(552,219)(556,219){9}
//: {10}(372,261)(372,219)(383,219){11}
//: {12}(173,261)(173,214)(183,214){13}
//: {14}(-69,261)(-69,219)(-38,219){15}
//: {16}(-170,265)(-170,213){17}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-195,285){13}
//: {14}(-199,285)(-237,285){15}
//: {16}(-197,287)(-197,347)(-167,347)(-167,336){17}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 8 10 7 -1 ]
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 11 0 ]
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  //: joint g54 (RegWrite) @(-170, 263) /w:[ 2 -1 1 16 ]
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 9 0 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 15 0 ]
  led g52 (.I(clk));   //: @(-167,329) /sn:0 /w:[ 17 ] /type:0
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 15 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 13 1 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 6 12 5 -1 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 4 14 3 -1 ]
  //: joint g55 (clk) @(-197, 285) /w:[ 13 -1 14 16 ]
  led g53 (.I(RegWrite));   //: @(-170,206) /sn:0 /w:[ 17 ] /type:0
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clk, clr, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Li0>clk(59/69) Li1>RegWr(47/69) Li2>SB[2:0](22/69) Li3>SA[2:0](11/69) Li4>SD[2:0](35/69) Ri0>clr(35/69) Bo0<BOUT[31:0](65/98) Bo1<AOUT[31:0](37/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module main;    //: root_module
supply0 w13;    //: /sn:0 {0}(45,134)(45,169){1}
supply0 w7;    //: /sn:0 {0}(157,281)(157,271)(172,271)(172,353)(219,353)(219,342){1}
supply0 [15:0] w20;    //: /sn:0 {0}(736,324)(694,324){1}
supply1 w12;    //: /sn:0 {0}(343,100)(343,142){1}
supply0 w32;    //: /sn:0 {0}(1340,241)(1340,214){1}
supply0 w35;    //: /sn:0 {0}(1033,-195)(1033,-150){1}
supply1 [15:0] w26;    //: /sn:0 /dp:1 {0}(682,354)(708,354)(708,344)(736,344){1}
supply0 [31:0] w9;    //: /sn:0 {0}(250,150)(329,150){1}
wire [31:0] w16;    //: /sn:0 {0}(1010,267)(917,267){1}
//: {2}(915,265)(915,-110)(1019,-110){3}
//: {4}(915,269)(915,297)(972,297)(972,318)(1002,318)(1002,356)(989,356){5}
wire [31:0] w6;    //: /sn:0 {0}(358,166)(495,166)(495,-142)(925,-142){1}
//: {2}(929,-142)(1019,-142){3}
//: {4}(927,-144)(927,-159)(1148,-159)(1148,-146)(1186,-146){5}
wire [31:0] w34;    //: /sn:0 /dp:1 {0}(1399,136)(1415,136)(1415,185){1}
//: {2}(1417,187)(1469,187){3}
//: {4}(1413,187)(1364,187){5}
wire [4:0] w25;    //: /sn:0 {0}(708,227)(737,227){1}
wire [5:0] w39;    //: /sn:0 {0}(921,365)(921,398)(1020,398)(1020,348)(1092,348){1}
wire [31:0] w36;    //: /sn:0 {0}(1215,-136)(1436,-136){1}
wire [5:0] w22;    //: /sn:0 /dp:1 {0}(635,114)(700,114)(700,21)(730,21)(730,6)(742,6){1}
wire w3;    //: /sn:0 {0}(4570,226)(4560,226){1}
wire [31:0] w0;    //: /sn:0 {0}(1186,189)(1296,189){1}
//: {2}(1300,189)(1329,189){3}
//: {4}(1298,191)(1298,224)(1388,224)(1388,207)(1469,207){5}
wire w30;    //: /sn:0 {0}(23964,4072)(23964,4082)(23954,4082){1}
wire [31:0] w29;    //: /sn:0 /dp:1 {0}(1112,166)(891,166){1}
wire w37;    //: /sn:0 {0}(552,175)(552,185)(563,185)(563,169)(588,169){1}
//: {2}(590,167)(590,-8)(742,-8){3}
//: {4}(590,171)(590,305)(695,305)(695,250){5}
wire w42;    //: /sn:0 {0}(982,-16)(1145,-16)(1145,-43)(1173,-43){1}
wire w18;    //: /sn:0 /dp:1 {0}(1346,87)(1346,70){1}
//: {2}(1348,68)(1391,68)(1391,131){3}
//: {4}(1346,66)(1346,57)(1347,57)(1347,44){5}
wire [3:0] w19;    //: /sn:0 {0}(1149,317)(1149,229){1}
wire [15:0] w23;    //: /sn:0 /dp:5 {0}(983,361)(921,361){1}
//: {2}(920,361)(794,361)(794,380)(752,380){3}
//: {4}(751,380)(647,380)(647,312)(635,312){5}
wire w10;    //: /sn:0 {0}(966,-31)(966,-78)(1452,-78)(1452,-123){1}
wire w54;    //: /sn:0 {0}(1194,-40)(1202,-40)(1202,-113){1}
wire w24;    //: /sn:0 {0}(752,375)(752,357){1}
wire [4:0] w21;    //: /sn:0 {0}(679,217)(661,217)(661,202){1}
//: {2}(661,198)(661,179)(716,179)(716,191)(737,191){3}
//: {4}(659,200)(635,200){5}
wire [4:0] w31;    //: /sn:0 {0}(679,237)(662,237)(662,236)(635,236){1}
wire [31:0] w1;    //: /sn:0 {0}(201,317)(173,317)(173,207)(73,207){1}
//: {2}(71,205)(71,182)(329,182){3}
//: {4}(69,207)(50,207){5}
wire w53;    //: /sn:0 /dp:1 {0}(1173,-38)(1161,-38)(1161,143){1}
wire w8;    //: /sn:0 {0}(343,201)(343,190){1}
wire w46;    //: /sn:0 {0}(18,118)(23,118)(23,120)(33,120){1}
//: {2}(35,118)(35,115){3}
//: {4}(35,122)(35,169){5}
wire w52;    //: /sn:0 /dp:1 {0}(874,118)(874,108)(919,108)(919,62){1}
wire [31:0] w44;    //: /sn:0 /dp:1 {0}(891,247)(942,247){1}
//: {2}(946,247)(1010,247){3}
//: {4}(944,245)(944,110)(1331,110)(1331,120)(1366,120)(1366,136)(1383,136){5}
wire [31:0] w27;    //: /sn:0 {0}(236,315)(631,315)(631,312){1}
//: {2}(631,311)(631,236){3}
//: {4}(631,235)(631,200){5}
//: {6}(631,199)(631,160){7}
//: {8}(631,159)(631,114){9}
//: {10}(631,113)(631,-174)(1305,-174)(1305,-156)(1436,-156){11}
wire [1:0] w17;    //: /sn:0 /dp:1 {0}(982,23)(1085,23)(1085,285)(1109,285)(1109,317){1}
wire [31:0] w28;    //: /sn:0 {0}(29,207)(-106,207)(-106,-218)(1507,-218)(1507,-146)(1465,-146){1}
wire w33;    //: /sn:0 {0}(1033,-102)(1033,-92){1}
wire w14;    //: /sn:0 {0}(-154,453)(38,453){1}
//: {2}(42,453)(847,453){3}
//: {4}(851,453)(1328,453)(1328,13)(1345,13)(1345,23){5}
//: {6}(849,451)(849,303){7}
//: {8}(40,451)(40,335){9}
wire w45;    //: /sn:0 /dp:1 {0}(1350,23)(1350,-25)(1161,-25)(1161,35)(982,35){1}
wire [15:0] w49;    //: /sn:0 /dp:1 {0}(765,334)(899,334)(899,351)(983,351){1}
wire [31:0] w41;    //: /sn:0 /dp:1 {0}(737,267)(553,267)(553,448)(1532,448)(1532,197)(1498,197){1}
wire w2;    //: /sn:0 {0}(1485,174)(1485,9)(982,9){1}
wire w48;    //: /sn:0 {0}(40,319)(40,245){1}
wire [31:0] w47;    //: /sn:0 /dp:1 {0}(1039,257)(1076,257)(1076,212)(1095,212)(1095,201)(1112,201){1}
wire [4:0] w15;    //: /sn:0 {0}(737,151)(682,151)(682,160)(635,160){1}
wire w55;    //: /sn:0 /dp:1 {0}(1346,103)(1346,161)(1347,161)(1347,164){1}
wire w38;    //: /sn:0 {0}(1026,234)(1026,47)(982,47){1}
wire w5;    //: /sn:0 {0}(-44,92)(-11,92){1}
//: {2}(-7,92)(806,92)(806,118){3}
//: {4}(-9,94)(-9,118)(2,118){5}
wire w43;    //: /sn:0 /dp:1 {0}(1427,245)(1442,245)(1442,229)(1428,229)(1428,44)(1445,44)(1445,-1)(982,-1){1}
wire [31:0] w40;    //: /sn:0 {0}(1048,-126)(1186,-126){1}
wire w51;    //: /sn:0 {0}(1411,245)(1381,245)(1381,261)(1354,261)(1354,214){1}
//: enddecls

  tran g44(.Z(w24), .I(w23[15]));   //: @(752,378) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:0
  register g4 (.Q(w1), .D(w28), .EN(w13), .CLR(w46), .CK(w48));   //: @(40,207) /sn:0 /R:1 /w:[ 5 0 1 5 1 ]
  //: joint g8 (w1) @(71, 207) /w:[ 1 2 4 -1 ]
  //: supply0 g47 (w20) @(688,324) /sn:0 /R:3 /w:[ 1 ]
  add g16 (.A(w16), .B(w6), .S(w40), .CI(w35), .CO(w33));   //: @(1035,-126) /sn:0 /R:1 /w:[ 3 3 0 1 0 ]
  tran g3(.Z(w31), .I(w27[15:11]));   //: @(629,236) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  //: joint g26 (w6) @(927, -142) /w:[ 2 4 1 -1 ]
  mux g17 (.I0(w6), .I1(w40), .S(w54), .Z(w36));   //: @(1202,-136) /sn:0 /R:1 /w:[ 5 1 1 0 ] /ss:0 /do:1
  add g2 (.A(w1), .B(w9), .S(w6), .CI(w12), .CO(w8));   //: @(345,166) /sn:0 /R:1 /w:[ 3 1 0 1 1 ]
  //: joint g30 (w0) @(1298, 189) /w:[ 2 -1 1 4 ]
  //: switch MEM_WRITE (w30) @(23964,4059) /R:3 /w:[ 0 ] /st:0
  tran g23(.Z(w22), .I(w27[31:26]));   //: @(629,114) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:1
  mux g39 (.I0(w44), .I1(w16), .S(w38), .Z(w47));   //: @(1026,257) /sn:0 /R:1 /w:[ 3 0 0 0 ] /ss:1 /do:1
  tran g1(.Z(w15), .I(w27[25:21]));   //: @(629,160) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  concat g24 (.I0(w23), .I1(w49), .Z(w16));   //: @(988,356) /sn:0 /w:[ 0 1 5 ] /dr:0
  mux g29 (.I0(w0), .I1(w34), .S(w2), .Z(w41));   //: @(1485,197) /sn:0 /R:1 /w:[ 5 3 0 1 ] /ss:1 /do:0
  not g60 (.I(w43), .Z(w51));   //: @(1421,245) /sn:0 /R:2 /w:[ 0 0 ]
  not g51 (.I(w14), .Z(w48));   //: @(40,329) /sn:0 /R:1 /w:[ 9 0 ]
  not g18 (.I(w5), .Z(w46));   //: @(8,118) /sn:0 /w:[ 5 0 ]
  mux g25 (.I0(w20), .I1(w26), .S(w24), .Z(w49));   //: @(752,334) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:1
  //: supply0 g10 (w7) @(157,287) /sn:0 /w:[ 0 ]
  //: joint g49 (w16) @(915, 267) /w:[ 1 2 -1 4 ]
  //: supply1 g6 (w12) @(354,100) /sn:0 /w:[ 0 ]
  not g50 (.I(w18), .Z(w55));   //: @(1346,93) /sn:0 /R:3 /w:[ 0 0 ]
  tran g9(.Z(w21), .I(w27[20:16]));   //: @(629,200) /sn:0 /R:2 /w:[ 5 5 6 ] /ss:1
  //: supply0 g7 (w9) @(244,150) /sn:0 /R:3 /w:[ 0 ]
  //: joint g68 (w46) @(35, 120) /w:[ -1 2 1 4 ]
  //: supply0 g31 (w32) @(1340,247) /sn:0 /w:[ 0 ]
  rom MemoRom (.A(w1), .D(w27), .OE(w7));   //: @(219,316) /sn:0 /w:[ 0 0 1 ] /mem:"/home/milax/Baixades/mult (1).mem"
  and g22 (.I0(w42), .I1(w53), .Z(w54));   //: @(1184,-40) /sn:0 /w:[ 1 0 0 ]
  //: joint g45 (w14) @(849, 453) /w:[ 4 6 3 -1 ]
  AC g41 (.AluOp(w17), .Funct(w39), .AluCtrl(w19));   //: @(1093, 318) /sz:(93, 70) /sn:0 /p:[ Ti0>1 Li0>1 To0<0 ]
  //: joint g54 (w14) @(40, 453) /w:[ 2 8 1 -1 ]
  UC g42 (.op(w22), .Jump(w10), .RegDst(w37), .RegWrite(w52), .AluSrc(w38), .MemWrite(w45), .AluOp(w17), .MemToReg(w2), .MemRead(w43), .Branch(w42));   //: @(743, -30) /sz:(238, 91) /sn:0 /p:[ Li0>1 To0<0 Lo0<3 Bo0<1 Ro0<1 Ro1<1 Ro2<0 Ro3<1 Ro4<1 Ro5<0 ]
  //: joint g40 (w34) @(1415, 187) /w:[ 2 1 4 -1 ]
  //: joint g69 (w5) @(-9, 92) /w:[ 2 -1 1 4 ]
  mux g12 (.I0(w21), .I1(w31), .S(w37), .Z(w25));   //: @(695,227) /sn:0 /R:1 /w:[ 0 0 5 0 ] /ss:0 /do:1
  and g28 (.I0(w45), .I1(w14), .Z(w18));   //: @(1347,34) /sn:0 /R:3 /w:[ 0 5 5 ]
  //: joint g46 (w44) @(944, 247) /w:[ 2 4 1 -1 ]
  tran g14(.Z(w23), .I(w27[15:0]));   //: @(629,312) /sn:0 /R:2 /w:[ 5 1 2 ] /ss:1
  //: switch g11 (w3) @(4588,226) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: supply0 g5 (w13) @(45,128) /sn:0 /R:2 /w:[ 0 ]
  clock g19 (.Z(w14));   //: @(-167,453) /sn:0 /w:[ 0 ] /omega:750 /phi:0 /duty:50
  //: joint g61 (w37) @(590, 169) /w:[ -1 2 1 4 ]
  tran g21(.Z(w39), .I(w23[5:0]));   //: @(921,359) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: supply0 g32 (w35) @(1033,-201) /sn:0 /R:2 /w:[ 0 ]
  mux g20 (.I0(w36), .I1(w27), .S(w10), .Z(w28));   //: @(1452,-146) /sn:0 /R:1 /w:[ 1 11 1 1 ] /ss:0 /do:0
  //: switch reset (w5) @(-61,92) /sn:0 /w:[ 0 ] /st:0
  //: joint g63 (w18) @(1346, 68) /w:[ 2 4 -1 1 ]
  ram g38 (.A(w0), .D(w34), .WE(w55), .OE(w51), .CS(w32));   //: @(1347,188) /sn:0 /w:[ 3 5 1 1 1 ]
  BRegs32x32 g0 (.RegWrite(w52), .clr(w5), .Read1(w15), .Read2(w21), .Write(w25), .WriteData(w41), .clk(w14), .Data1(w29), .Data2(w44));   //: @(738, 119) /sz:(152, 183) /sn:0 /p:[ Ti0>0 Ti1>3 Li0>0 Li1>3 Li2>1 Li3>0 Bi0>7 Ro0<1 Ro1<0 ]
  ALU g15 (.B(w47), .A(w29), .ALU_C(w19), .Z(w53), .S(w0));   //: @(1113, 144) /sz:(72, 84) /sn:0 /p:[ Li0>1 Li1>0 Bi0>1 To0<1 Ro0<0 ]
  //: supply1 g48 (w26) @(682,343) /sn:0 /R:1 /w:[ 0 ]
  led g62 (.I(w37));   //: @(552,168) /sn:0 /w:[ 0 ] /type:0
  bufif1 g37 (.Z(w34), .I(w44), .E(w18));   //: @(1389,136) /sn:0 /w:[ 0 5 3 ]
  //: joint g13 (w21) @(661, 200) /w:[ -1 2 4 1 ]

endmodule
